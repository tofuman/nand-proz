module steuerwerk(control, status, instructionbus);
