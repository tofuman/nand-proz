module memman (addruper, addrlower, word)

